
module calculator_final (
	clk_clk,
	output_all_external_connection_export,
	input_6_external_connection_export,
	input_5_external_connection_export,
	input_4_external_connection_export,
	input_3_external_connection_export,
	input_2_external_connection_export,
	input_1_external_connection_export);	

	input		clk_clk;
	output	[7:0]	output_all_external_connection_export;
	input		input_6_external_connection_export;
	input		input_5_external_connection_export;
	input		input_4_external_connection_export;
	input		input_3_external_connection_export;
	input	[3:0]	input_2_external_connection_export;
	input	[3:0]	input_1_external_connection_export;
endmodule

module bin2bcd(clk1,tens,ones,
    bin
    );

    input clk1;
	 output[3:0] tens;
	 output[3:0] ones;
    //input ports and their sizes
    input [7:0] bin;
    //output ports and, their size
    reg [11:0] bcd;
    //Internal variables 
     reg [3:0] i;   
     
     //Always block - implement the Double Dabble algorithm
     always @(posedge clk1)
        begin
            bcd = 0; //initialize bcd to zero.
            for (i = 0; i < 8; i = i+1) //run for 8 iterations
            begin
                bcd = {bcd[10:0],bin[7-i]}; //concatenation
                    
                //if a hex digit of 'bcd' is more than 4, add 3 to it.  
                if(i < 7 && bcd[3:0] > 4) 
                    bcd[3:0] = bcd[3:0] + 3;
                if(i < 7 && bcd[7:4] > 4)
                    bcd[7:4] = bcd[7:4] + 3;
                if(i < 7 && bcd[11:8] > 4)
                    bcd[11:8] = bcd[11:8] + 3;  
            end
        end     
		  assign tens[3:0] = bcd[7:4];
		  assign ones[3:0] = bcd[3:0];
             
endmodule 